`timescale 1ns/1ns

module TEST1;

reg [3:0] a,b;
reg k;
wire [8:0] cout;
subBCD T_1(a,b,k,cout);
initial begin

a=4'b0000; b=4'b0000; k=0;
#10 a=4'b0001; b=4'b0001; k=0; //1+1
#10 a=4'b0011; b=4'b0001; k=0;//3+1
#10 a=4'b0111; b=4'b0001; k=0;//7+1
#10 a=4'b1111; b=4'b0001; k=0;//-1+1
#10 a=4'b0111; b=4'b0111; k=0;//7+7
#10 a=4'b0000; b=4'b0001; k=1;//0-1
#10 a=4'b0111; b=4'b0111; k=1;//7-7
#10 a=4'b1001; b=4'b0111; k=1;//-7-7
#10 a=4'b1001; b=4'b0001; k=1;//-7-1
#10 a=4'b0111; b=4'b1000; k=1;//7-8
#10 $finish;
end
endmodule
